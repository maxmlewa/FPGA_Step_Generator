`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Module Name: step_counter
// Project Name: Step Generator
// Target Devices: Basys 3 (Artix 7)
// Description: Counter triggered by a clean pulse input. Counts from 0 to steps -1.
//              Wraps around to 0. Freezes at 0 if steps = 0
// 
// Dependencies: None
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments: Couner resets on rising edge of rst input.
// 
//////////////////////////////////////////////////////////////////////////////////


module step_counter(

    );
endmodule
