`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Module Name: step_selector
// Project Name: Step Generator
// Target Devices: XXXX
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module step_selector(

    );
endmodule
