`timescale 1ns / 1ps
////////////////////////////////////////////////////////////////////////////////// 
// Module Name: testbench_step_selector
// Project Name: Step Generator
// Target Devices: Basys 3 (Artix 7)
// Description: Verifies correct priority encoding of the 10-bit switch input.
//              Tests single active inputs and multiple simultaneous inputs,
//              and no input case. Outputs should reflect the highest active bit
// 
// Dependencies: step_selector.v
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//  - All switches tested from highest to lowest priority.
//  - Multi-active input test ensures correcct priority encoding.
//  - Zero-input condition verified
// 
//////////////////////////////////////////////////////////////////////////////////


module testbench_step_selector(

    );
endmodule
