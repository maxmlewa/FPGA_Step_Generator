`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Module Name: step_selector
// Project Name: Step Generator
// Target Devices: Basys 3 (Artix 7)
// Description: Encodes active switch input (SW[9:0]) into a 4-bit number (range 1-10)
//              using priority encoding logic, with descending priority
// 
// Dependencies: None
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments: If no switches are active, outputs 0.
// 
//////////////////////////////////////////////////////////////////////////////////


module step_selector(

    );
endmodule
