`timescale 1ns / 1ps
////////////////////////////////////////////////////////////////////////////////// 
// Module Name: top_module_step_gen
// Project Name: Step Generator
// Target Devices: XXXX
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module top_module_step_gen(

    );
endmodule
