`timescale 1ns / 1ps
////////////////////////////////////////////////////////////////////////////////// 
// Module Name: top_module_step_gen
// Project Name: Step Generator
// Target Devices: Basys 3 (Artix 7)
// Description: Integrates all the modules to implement the step generator triggered
//              by an external clock signal. Output binary step count and displays the
//              step configuration.
// 
// Dependencies: step_selector, step_counter, edge_detector_debounced, seven_seg_display
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments: The counter output will be routed to an external DAC
// 
//////////////////////////////////////////////////////////////////////////////////


module top_module_step_gen(

    );
endmodule
