`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Module Name: step_counter
// Project Name: Step Generator
// Target Devices: XXXX
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module step_counter(

    );
endmodule
