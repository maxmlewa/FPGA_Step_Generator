`timescale 1ns / 1ps
////////////////////////////////////////////////////////////////////////////////// 
// Module Name: seven_seg_display
// Project Name: Step Generator
// Target Devices: Basys 3 (Artix 7)
// Description: Displays the current step configuration (1-10) on the rightmost
//              7-segment digit (an[0]). Supports digits 0-9 and 10 ("A").
// 
// Dependencies: None
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments: Display is active-low. Only an[0] is enabled.
// 
//////////////////////////////////////////////////////////////////////////////////


module seven_seg_display(

    );
endmodule
