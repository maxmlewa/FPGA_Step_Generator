`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Module Name: testbench_seven_seg_display
// Project Name: Step Generator
// Target Devices: Basys 3 (Atrix 7)
// Tool Versions: Vivado 2025
// Description: Verifies that each input maps to the LED pattern correctly
//              Ensure that inactive or  undefined values are disabled
// 
// Dependencies: seven_seg_display.v
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// - Segment outputs areactive-low
// - Rightmost display digit (an[0])is active, others off
//////////////////////////////////////////////////////////////////////////////////


module testbench_seven_seg_display(

    );
endmodule
